library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity dram_controller is port(
);
end dram_controller;

architecture dram_controller_arch of dram_controller is
begin
end architecture;