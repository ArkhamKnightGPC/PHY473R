library ieee;

use ieee.std_logic_1164.all;

entity camera_controller is port(
);
end camera_controller;

architecture camera_controller_arch of camera_controller is
begin
end architecture;